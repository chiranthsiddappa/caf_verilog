`timescale 1ns/1ns

module reference_buffer #(parameter buffer_length = 10,
                          parameter buffer_bits = 4,
                          parameter i_bits = 12,
                          parameter q_bits = 12
                          )
   (input clk,
    input                            m_axis_tready,
    input                            m_axis_index_tvalid,
    input [buffer_bits - 1:0]        m_axis_index_tdata,
    output reg                       s_axis_data_tready,
    output reg signed [i_bits - 1:0] i,
    output reg signed [q_bits - 1:0] q,
    output reg                       s_axis_data_tvalid
    );

   reg                               m_valid;
   reg [i_bits + q_bits - 1:0]       buffer [0:buffer_length - 1];
   reg [buffer_bits - 1:0]           addr_buffer;

   initial begin
      $readmemb("{{ reference_buffer_filename }}", buffer);
      s_axis_data_tvalid = 1'b0;
      s_axis_data_tready = 1'b1;
      m_valid = 1'b0;
   end

   always @(posedge clk) begin
      m_valid <= m_axis_index_tvalid & m_axis_tready;
      addr_buffer <= m_axis_index_tdata;
   end

   always @(posedge clk) begin
      if (m_valid && (addr_buffer < buffer_length)) begin
         i <= buffer[addr_buffer] >> q_bits;
         q <= buffer[addr_buffer] & ((1'b1 << q_bits) - 1);
         s_axis_data_tvalid <= 1'b1;
      end else begin
         s_axis_data_tvalid <= 1'b0;
      end
   end
endmodule // reference_buffer
